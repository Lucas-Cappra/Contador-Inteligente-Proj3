LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY SOMADOR_BCD_12 IS
	PORT(
	A_BCD_U, B_BCD_STEP: IN STD_LOGIC_VECTOR(3 DOWNTO 0); --A � O NUMEROMAX/MIN B VAI SER O STE
	A_BCD_D, B_BCD_D: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	A_BCD_C, B_BCD_C: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	CI_BCD: IN STD_LOGIC;
	CO_BCD: OUT STD_LOGIC;
	S_BCD_U: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	S_BCD_D: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	S_BCD_C: OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
);
END SOMADOR_BCD_12;

ARCHITECTURE SOMA_12BITS_BCD OF SOMADOR_BCD_12 IS
	COMPONENT Somador_BCD IS
		PORT(
        	A, B: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        	CI: IN STD_LOGIC;
        	S: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
        	CO: OUT STD_LOGIC
    	);
	END COMPONENT;
	
	SIGNAL CO_1, CO_2: STD_LOGIC;
BEGIN

SS_12_U : Somador_BCD PORT MAP(A_BCD_U, B_BCD_STEP, '0', S_BCD_U, CO_1);
SS_12_D : Somador_BCD PORT MAP(A_BCD_D, "0000", CO_1,   S_BCD_D, CO_2);
SS_12_C : Somador_BCD PORT MAP(A_BCD_C, "0000", CO_2,   S_BCD_C, CO_BCD);


END ARCHITECTURE;