LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY SUBTRATOR IS
	PORT(
	A_BCD_U, B_BCD_STEP: IN STD_LOGIC_VECTOR(3 DOWNTO 0); --A � O NUMEROMAX/MIN B VAI SER O STE
	A_BCD_D: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	A_BCD_C: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	CI_BCD: IN STD_LOGIC;
	CO_BCD: OUT STD_LOGIC;
	S_BCD_U: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	S_BCD_D: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	S_BCD_C: OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
);
END SUBTRATOR;

ARCHITECTURE SUB_12_P OF SUBTRATOR IS
	COMPONENT SUB_BCD_COMP IS
	PORT(
	A, B: IN STD_LOGIC_VECTOR(3 DOWNTO 0); -- A SAIDA REG MAX/MIN E B VAI SER O STEP
	CI: IN STD_LOGIC;
	SINAL: OUT STD_LOGIC;
	S: OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
);
	END COMPONENT;
	
	SIGNAL CO_1, CO_2: STD_LOGIC;
BEGIN

SS_12_U : SUB_BCD_COMP PORT MAP(A_BCD_U, B_BCD_STEP, '0',CO_1, S_BCD_U);
SS_12_D : SUB_BCD_COMP PORT MAP(A_BCD_D, "0000", CO_1, CO_2,S_BCD_D);
SS_12_C : SUB_BCD_COMP PORT MAP(A_BCD_C, "0000", CO_2, CO_BCD, S_BCD_C);

END ARCHITECTURE;
