LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY SUBTRATOR_BCD_12 IS
    PORT(
    A_BCD_U, B_BCD_STEP: IN STD_LOGIC_VECTOR(3 DOWNTO 0); --A � O NUMEROMAX/MIN B VAI SER O STE
    A_BCD_D: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    A_BCD_C: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    CO_BCD: OUT STD_LOGIC;
    S_BCD_U: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    S_BCD_D: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    S_BCD_C: OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
);
END SUBTRATOR_BCD_12;

ARCHITECTURE SUB_12BITS_BCD OF SUBTRATOR_BCD_12 IS
	COMPONENT SUB_BCD_COMP IS
		PORT(
		A, B: IN STD_LOGIC_VECTOR(3 DOWNTO 0); -- A SAIDA REG MAX/MIN E B VAI SER O STEP
		CI: IN STD_LOGIC;
		SINAL: OUT STD_LOGIC;
		S: OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);

	END COMPONENT;


	COMPONENT Somador_4Bits IS
		Port(
        	A_S4, B_S4: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        	CI_S4: IN STD_LOGIC;
        	S_S4: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
        	CO_S4: OUT STD_LOGIC
     	);
    	END COMPONENT;

    SIGNAL CO_1, CO_2, CO_BCD_AUX: STD_LOGIC;
    SIGNAL CO_1_AUX, CO_2_AUX: STD_LOGIC_VECTOR(3 DOWNTO 0);
    SIGNAL S_BCD_U_AUX, S_BCD_D_AUX, S_BCD_C_AUX: STD_LOGIC_VECTOR(3 DOWNTO 0);
    SIGNAL S_BCD_U1, S_BCD_U1_RES: STD_LOGIC_VECTOR(3 DOWNTO 0);
    SIGNAL S_BCD_D2, S_BCD_D2_RES: STD_LOGIC_VECTOR(3 DOWNTO 0);
    SIGNAL S_BCD_C3, S_BCD_C3_RES: STD_LOGIC_VECTOR(3 DOWNTO 0);
    SIGNAL C0_AUX1: STD_LOGIC_VECTOR(5 DOWNTO 0);
    SIGNAL SOMA1, SOMA2, SOMA3, SOMAR1, SOMAR2, SOMAR3: STD_LOGIC_VECTOR(3 DOWNTO 0);
    
BEGIN

--UNIDADE
SS_12_U : SUB_BCD_COMP PORT MAP(A_BCD_U, B_BCD_STEP, '0', CO_1, S_BCD_U_AUX);

--S_BCD_U <= NOT(CO_1) AND S_BCD_U_AUX; --SE CO_1 = '0', RECEBE O VALOR NORMAL DA SA�DA
--COMPLEMENTO A 2 QUANDO NUMERO � NEGATIVO E SOMA 10
S_BCD_U1(3) <= CO_1 XOR S_BCD_U_AUX(3);
S_BCD_U1(2) <= CO_1 XOR S_BCD_U_AUX(2);
S_BCD_U1(1) <= CO_1 XOR S_BCD_U_AUX(1);
S_BCD_U1(0) <= CO_1 XOR S_BCD_U_AUX(0);

SOMAR1(3) <= '0';
SOMAR1(2) <= '0';
SOMAR1(1) <= '0';
SOMAR1(0) <= '1' AND CO_1;

AUX1: Somador_4Bits PORT MAP (S_BCD_U1, SOMAR1, '0', S_BCD_U1_RES, C0_AUX1(5));

SOMA1(3) <= '1' AND CO_1;
SOMA1(2) <= '0';
SOMA1(1) <= '1' AND CO_1;
SOMA1(0) <= '0';

AUX2 : Somador_4Bits PORT MAP (S_BCD_U1_RES, SOMA1, '0', S_BCD_U, C0_AUX1(4));

--DEZENA
CO_1_AUX(3) <= '0';
CO_1_AUX(2) <= '0';
CO_1_AUX(1) <= '0';
CO_1_AUX(0) <= CO_1 AND '1';
SS_12_D : SUB_BCD_COMP PORT MAP(A_BCD_D, CO_1_AUX, CO_1, CO_2, S_BCD_D_AUX);

--COMPLEMENTO A 2 QUANDO NUMERO � NEGATIVO E SOMA 10
S_BCD_D2(3) <= CO_2 XOR S_BCD_D_AUX(3);
S_BCD_D2(2) <= CO_2 XOR S_BCD_D_AUX(2);
S_BCD_D2(1) <= CO_2 XOR S_BCD_D_AUX(1);
S_BCD_D2(0) <= CO_2 XOR S_BCD_D_AUX(0);

SOMAR2(3) <= '0';
SOMAR2(2) <= '0';
SOMAR2(1) <= '0';
SOMAR2(0) <= '1' AND CO_2;

AUX3: Somador_4Bits PORT MAP (S_BCD_D2, SOMAR2, '0', S_BCD_D2_RES, C0_AUX1(3));

SOMA2(3) <= '1' AND CO_2;
SOMA2(2) <= '0';
SOMA2(1) <= '1' AND CO_2;
SOMA2(0) <= '0';

AUX4 : Somador_4Bits PORT MAP (S_BCD_D2_RES, SOMA2, '0', S_BCD_D, C0_AUX1(2));

--CENTENA
CO_2_AUX(3) <= '0';
CO_2_AUX(2) <= '0';
CO_2_AUX(1) <= '0';
CO_2_AUX(0) <= CO_2 AND '1';
SS_12_C : SUB_BCD_COMP PORT MAP(A_BCD_C, CO_2_AUX, CO_2,   CO_BCD_AUX, S_BCD_C);
END ARCHITECTURE;
