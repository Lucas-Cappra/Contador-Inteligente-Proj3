LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY SUBTRATOR_COMPLETO_12Bits IS
    PORT(
        A_U, BCD_STEP: IN STD_LOGIC_VECTOR(3 DOWNTO 0); -- A � O NUMEROMAX/MIN B VAI SER O STE
        A_D: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        A_C: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	CO_D: OUT STD_LOGIC;
        S_U: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
        S_D: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
        S_C: OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
    );
END SUBTRATOR_COMPLETO_12Bits;

ARCHITECTURE SUBTRATOR_COMPLETO_12Bits OF SUBTRATOR_COMPLETO_12Bits IS
    COMPONENT SUBTRATOR IS -- A_U> STEP
	PORT(
	A_BCD_U, B_BCD_STEP: IN STD_LOGIC_VECTOR(3 DOWNTO 0); --A � O NUMEROMAX/MIN B VAI SER O STE
	A_BCD_D: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	A_BCD_C: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	CI_BCD: IN STD_LOGIC;
	CO_BCD: OUT STD_LOGIC;
	S_BCD_U: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	S_BCD_D: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	S_BCD_C: OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
);
    END COMPONENT;

    COMPONENT SUBTRATOR_BCD_12 IS -- STEP> A_U
    PORT(
    A_BCD_U, A_BCD_D, A_BCD_C: IN STD_LOGIC_VECTOR(3 DOWNTO 0); --A � O NUMEROMAX/MIN B VAI SER O STE
    B_BCD_STEP: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    S_BCD_U: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    S_BCD_D: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    S_BCD_C: OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
);
    END COMPONENT;

    COMPONENT MUX_4X1_4BITS IS
	PORT (
        A, B : in  STD_LOGIC_VECTOR(3 DOWNTO 0);
        C    : in  STD_LOGIC;
        Y    : out STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
    END COMPONENT;

    SIGNAL A_MAIOR_STEP: STD_LOGIC; 
    SIGNAL S_U_AUX, S_D_AUX, S_C_AUX: STD_LOGIC_VECTOR (3 DOWNTO 0); --U1 VAI SER A_U>STEP E U2 VAI SER STEP> A_U
    SIGNAL S_U_AUX_2, S_C_AUX_2, S_D_AUX_2: STD_LOGIC_VECTOR (3 DOWNTO 0);
    SIGNAL S_Y_U, S_Y_D, S_Y_C: STD_LOGIC_VECTOR (3 DOWNTO 0);
    
BEGIN

A_U1: SUBTRATOR_BCD_12 PORT MAP (A_U, BCD_STEP, A_D, A_C, S_U_AUX, S_D_AUX, S_C_AUX);
A_U2: SUBTRATOR PORT MAP (A_U, BCD_STEP, A_D, A_C, '0', CO_D ,S_U_AUX_2, S_D_AUX_2, S_C_AUX_2);


A_MAIOR_STEP <= ((not(A_U(3)) and BCD_STEP(3)) or 
 		((A_U(3) xnor BCD_STEP(3)) and not(A_U(2)) and BCD_STEP(2)) or 
        	((A_U(3) xnor BCD_STEP(3)) and (A_U(2) xnor BCD_STEP(2)) and  not(A_U(1)) and BCD_STEP(1)) or 
        	((A_U(3) xnor BCD_STEP(3)) and (A_U(2) xnor BCD_STEP(2)) and  (A_U(1) xnor BCD_STEP(1)) and  not(A_U(0))�and�BCD_STEP(0)));

MUX_U: MUX_4X1_4BITS PORT MAP(S_U_AUX, S_U_AUX_2, A_MAIOR_STEP, S_Y_U);
MUX_D: MUX_4X1_4BITS PORT MAP(S_D_AUX, S_D_AUX_2, A_MAIOR_STEP, S_Y_D);
MUX_C: MUX_4X1_4BITS PORT MAP(S_C_AUX, S_C_AUX_2, A_MAIOR_STEP, S_Y_C);

S_U <= S_Y_U;
S_D <= S_Y_D;
S_C <= S_Y_C;

END ARCHITECTURE;