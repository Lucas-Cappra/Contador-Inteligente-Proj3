LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY SUB_BCD_COMP IS
	PORT(
	A, B: IN STD_LOGIC_VECTOR(3 DOWNTO 0); -- A SAIDA REG MAX/MIN E B VAI SER O STEP
	CI: IN STD_LOGIC;
	SINAL: OUT STD_LOGIC;
	S: OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
);

END SUB_BCD_COMP;

ARCHITECTURE SUB_BCD OF SUB_BCD_COMP IS

COMPONENT Somador_4Bits IS
    Port(
        A_S4, B_S4: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        CI_S4: IN STD_LOGIC;
        S_S4: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
        CO_S4: OUT STD_LOGIC
    );
END COMPONENT;

SIGNAL B_XOR: STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL COS4_1, COS4_2, COS4_3, COS4_4: STD_lOGIC; -- CARRY OUT DE SAIDA DOS SOMADORES DE 4 BITS
SIGNAL S4_1, S4_2, S4_3, S4_4_AUX: STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL ES4_3, ES4_4: STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL CI_S4_AUX: STD_LOGIC;

BEGIN

B_XOR <= B XOR "1111";

I1 : Somador_4bits PORT MAP ("1010", B_XOR, '0', S4_1, COS4_1);
COS4_1 <= '0';


I2: Somador_4bits PORT MAP (A, S4_1, '0', S4_2, COS4_2);

--CONFIGURACAO NA SAIDA DO SOMADOR 2 COM O CARRY OUT
ES4_3(3) <= '0';
ES4_3(2) <= (S4_2(1) AND S4_2(3)) OR (S4_2(2) AND S4_2(3)) OR COS4_2;
ES4_3(1) <= (S4_2(1) AND S4_2(3)) OR (S4_2(2) AND S4_2(3)) OR COS4_2;
ES4_3(0) <= '0';


--CONFIGURACAO ENTRADA SOMADOR 4
ES4_4(3) <= NOT((S4_2(1) AND S4_2(3)) OR (S4_2(2) AND S4_2(3)) OR COS4_2);
ES4_4(2) <= '0';
ES4_4(1) <= NOT((S4_2(1) AND S4_2(3)) OR (S4_2(2) AND S4_2(3)) OR COS4_2);
ES4_4(0) <= '0'; 

S4_4_AUX(3) <= S4_3(3) XOR NOT((S4_2(1) AND S4_2(3)) OR (S4_2(2) AND S4_2(3)) OR COS4_2);
S4_4_AUX(2) <= S4_3(2) XOR NOT((S4_2(1) AND S4_2(3)) OR (S4_2(2) AND S4_2(3)) OR COS4_2);
S4_4_AUX(1) <= S4_3(1) XOR NOT((S4_2(1) AND S4_2(3)) OR (S4_2(2) AND S4_2(3)) OR COS4_2);
S4_4_AUX(0) <= S4_3(0) XOR NOT((S4_2(1) AND S4_2(3)) OR (S4_2(2) AND S4_2(3)) OR COS4_2);

CI_S4_AUX <= (S4_2(1) AND S4_2(3)) OR (S4_2(2) AND S4_2(3)) OR COS4_2;

--VOLTA A REALIZAR AS SOMAS
I3: Somador_4bits PORT MAP(ES4_3, S4_2, '0', S4_3, COS4_3);
COS4_3 <= '0';

I4: Somador_4bits PORT MAP(ES4_4, S4_4_AUX, CI_S4_AUX, S, COS4_4);

--SINAL DO NUMERO NA SAIDA DO SUBTRATOR
SINAL <= NOT((S4_2(1) AND S4_2(3)) OR (S4_2(2) AND S4_2(3)) OR COS4_2);

END ARCHITECTURE;
